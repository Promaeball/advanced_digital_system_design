* nand.cir

.subckt nand a b out vdd vss params: tplv=1 tpwv=1 tnlv=1 tnwv=1 tpotv=1 tnotv=1
M1 vdd a out vdd tp L={tplv * 65n} W={tpwv * 160n} 
+ AS=75.3f AD=75.3f PS=1.23u PD=1.23u
M2 vdd b out vdd tp L={tplv * 65n} W={tpwv * 185n} 
+ AS=75.3f AD=75.3f PS=1.23u PD=1.23u
M3 out a c c tn L={tnlv * 65n} W={tnwv * 130n} 
+ AS=75.3f AD=75.3f PS=1.12u PD=1.23u
M4 c b vss vss tn L={tnlv * 65n} W={tnwv * 130n} 
+ AS=75.3f AD=75.3f PS=1.12u PD=1.23u

.model tp pmos level=54 version=4.8.2 TOXE={tpotv * 1.95n}
.model tn nmos level=54 version=4.8.2 TOXE={tnotv * 1.85n}

.ends nand