* inverter

.subckt inverter in out vdd vss params: tplv=1 tpwv=1 tnlv=1 tnwv=1 tpotv=1 tnotv=1
M1 vdd in out vdd tp L={tplv * 65n} W={tpwv * 220n} 
+ AS=75.3f AD=75.3f PS=1.23u PD=1.23u
M2 out in vss vss tn L={tnlv * 65n} W={tnwv * 130n} 
+ AS=75.3f AD=75.3f PS=1.12u PD=1.23u

.model tp pmos level=54 version=4.8.2 TOX={tpotv * 1.95n}
.model tn nmos level=54 version=4.8.2 TOX={tnotv * 1.85n}

.ends inverter
