*ring_oscillator_6
.include nand.cir
.include inverter.cir
.subckt ring_oscillator_6 enable output vdd vss
X1 enable output n0 vdd vss nand tplv=1.076802 tpwv=0.989002 tnln=1.074132 tnwn=0.984710 tpotv=0.919926 tnotv=1.023770
X2 n0 n1 vdd vss inverter tplv=1.012438 tpwv=0.928178 tnln=0.977783 tnwn=0.944035 tpotv=1.013361 tnotv=0.921488
X3 n1 n2 vdd vss inverter tplv=0.982427 tpwv=0.976635 tnln=0.973989 tnwn=1.014305 tpotv=1.015101 tnotv=0.931186
X4 n2 n3 vdd vss inverter tplv=0.951478 tpwv=1.007650 tnln=0.964428 tnwn=0.924112 tpotv=0.974615 tnotv=0.986384
X5 n3 n4 vdd vss inverter tplv=1.007139 tpwv=1.042231 tnln=0.943260 tnwn=0.953883 tpotv=1.040426 tnotv=0.998159
X6 n4 n5 vdd vss inverter tplv=1.071122 tpwv=0.981979 tnln=1.053438 tnwn=0.928719 tpotv=1.046592 tnotv=0.985211
X7 n5 n6 vdd vss inverter tplv=1.094084 tpwv=1.029505 tnln=1.018775 tnwn=0.982010 tpotv=0.913047 tnotv=1.007262
X8 n6 n7 vdd vss inverter tplv=1.003001 tpwv=0.989870 tnln=0.970669 tnwn=0.877433 tpotv=1.026259 tnotv=1.032558
X9 n7 n8 vdd vss inverter tplv=1.038563 tpwv=0.996270 tnln=0.994389 tnwn=1.031855 tpotv=1.000429 tnotv=0.936839
X10 n8 n9 vdd vss inverter tplv=1.022602 tpwv=1.036603 tnln=0.985405 tnwn=0.998260 tpotv=1.008177 tnotv=0.983085
X11 n9 n10 vdd vss inverter tplv=0.953515 tpwv=0.963984 tnln=0.888779 tnwn=1.068965 tpotv=1.001183 tnotv=0.944279
X12 n10 n11 vdd vss inverter tplv=0.991272 tpwv=0.931251 tnln=1.026005 tnwn=0.979879 tpotv=1.084124 tnotv=0.980917
X13 n11 output vdd vss inverter tplv=0.983323 tpwv=0.991010 tnln=1.091388 tnwn=1.007820 tpotv=0.979483 tnotv=0.965705
.ends ring_oscillator_6
