* NAND gate using BSIM4
* File name nand.cir

* Voltage Supply
VDD VDD 0 1.0V

* Inputs
Vin1 IN1 0 PULSE (0 1.0 0 1n 1n 5n 10n) * Input pulse 1
Vin2 IN2 0 PULSE (0 1.0 0 1n 1n 5n 10n) * Input pulse 2

* Output Load
CL OUT 0 1f        

* Transistor Parameters
.model tn nmos BSIM4 level=54 version=4.8.2
.model tp pmos BSIM4 level=54 version=4.8.2

* NMOS Transistors
M1 OUT IN1 N1 0 NMOS W=130n L=50n
M2 OUT IN2 N1 0 NMOS W=130n L=50n

* PMOS Transistors
M3 OUT IN1 VDD VDD PMOS W=260n L=50n
M4 OUT IN2 VDD VDD PMOS W=260n L=50n
