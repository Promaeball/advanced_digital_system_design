*ring_oscillator_2
.include nand.cir
.include inverter.cir
.subckt ring_oscillator_2 enable output vdd vss
X1 enable output n0 vdd vss nand tplv=0.948158 tpwv=1.061308 tnln=0.895019 tnwn=1.009856 tpotv=0.961972 tnotv=1.038562
X2 n0 n1 vdd vss inverter tplv=0.950490 tpwv=1.009969 tnln=1.044809 tnwn=0.944979 tpotv=1.006718 tnotv=1.059439
X3 n1 n2 vdd vss inverter tplv=0.966296 tpwv=1.064987 tnln=1.044805 tnwn=0.913158 tpotv=1.035398 tnotv=1.093812
X4 n2 n3 vdd vss inverter tplv=1.055355 tpwv=1.021487 tnln=1.087745 tnwn=1.012733 tpotv=1.009596 tnotv=1.023991
X5 n3 n4 vdd vss inverter tplv=0.968482 tpwv=1.066314 tnln=1.036503 tnwn=0.974149 tpotv=0.966198 tnotv=1.074252
X6 n4 n5 vdd vss inverter tplv=1.063938 tpwv=0.950674 tnln=0.952756 tnwn=0.958307 tpotv=0.920428 tnotv=1.032471
X7 n5 n6 vdd vss inverter tplv=0.984925 tpwv=1.072294 tnln=0.993054 tnwn=1.059687 tpotv=0.953817 tnotv=0.997344
X8 n6 n7 vdd vss inverter tplv=1.078278 tpwv=0.979210 tnln=1.009659 tnwn=1.035276 tpotv=1.015727 tnotv=0.960054
X9 n7 n8 vdd vss inverter tplv=1.076576 tpwv=0.939143 tnln=1.039959 tnwn=0.937453 tpotv=0.954494 tnotv=0.948815
X10 n8 n9 vdd vss inverter tplv=1.014174 tpwv=0.857283 tnln=1.037809 tnwn=0.920402 tpotv=1.034520 tnotv=1.030751
X11 n9 n10 vdd vss inverter tplv=1.054037 tpwv=1.083032 tnln=1.016012 tnwn=0.949014 tpotv=1.029710 tnotv=0.998442
X12 n10 n11 vdd vss inverter tplv=0.977529 tpwv=1.060613 tnln=1.008170 tnwn=0.993138 tpotv=0.919535 tnotv=1.028127
X13 n11 output vdd vss inverter tplv=0.969867 tpwv=1.084281 tnln=0.992791 tnwn=0.998442 tpotv=1.053872 tnotv=1.006279
.ends ring_oscillator_2
