* NAND gate using BSIM4
* File name nand.cir

* Voltage Supply
VDD VDD 0 1.0V

* Inputs
Vin1 IN1 0 PULSE (0 1.0 0 1n 1n 5n 10n) * Input pulse 1
Vin2 IN2 0 PULSE (0 1.0 0 1n 1n 5n 10n) * Input pulse 2

* Output Load
CL OUT 0 1f        

* Transistor Parameters
.model tn nmos level=54 version=4.8.2 TOX=1.85n
.model tp pmos level=54 version=4.8.2 TOX=1.95n

* PMOS
M1 out in vdd vdd tp L=50n W=260n
+ AS=75.3f AD=75.3f PS=1.23u PD=1.23u
M2 out in vdd vdd tp L=50n W=260n
+ AS=75.3f AD=75.3f PS=1.23u PD=1.23u

* NMOS
M3 out in vss vss tn L=50n W=260n
+ AS=75.3f AD=75.3f PS=1.12u PD=1.23u
M4 out in vss vss tn L=50n W=260n
+ AS=75.3f AD=75.3f PS=1.12u PD=1.23u
