* Inverter with Parameters
.subckt inverter in out vdd vss L_pmos=65n W_pmos=130n L_nmos=65n W_nmos=130n TOX_pmos=1.95n TOX_nmos=1.85n

M1 out in vdd vdd tp L={L_pmos} W={W_pmos}
+ AS=75.3f AD=75.3f PS=1.23u PD=1.23u

M2 out in vss vss tn L={L_nmos} W={W_nmos}
+ AS=75.3f AD=75.3f PS=1.12u PD=1.23u

* BSIM4 4.8.2 models
.model tp PMOS level=54 version=4.8.2 TOX={TOX_pmos}
.model tn NMOS level=54 version=4.8.2 TOX={TOX_nmos}
.ends inverter
