* Inverter Model with BSIM4 and Parametric Variations
* Define process variation parameters
.param tplv=0.18u          * PMOS transistor length variation
.param tpwv=1.0u           * PMOS transistor width variation
.param tnln=0.18u          * NMOS transistor length variation
.param tnwn=1.0u           * NMOS transistor width variation
.param tpotv=2.0e-9        * PMOS transistor oxide thickness variation
.param tnotv=2.0e-9        * NMOS transistor oxide thickness variation

* Power Supply
VDD vdd 0 1.8V

* Input Signal
Vin in 0 PULSE(0 1.8 0 1n 1n 5n 10n)

* NMOS Transistor (BSIM4 Model)
M1 out in 0 0 NMOS L='tnln+tplv' W='tnwn+tpwv'
.model NMOS nmos level=54
+ toxe=tnotv                * NMOS transistor oxide thickness variation
+ ...                       * Additional NMOS BSIM4 parameters as needed

* PMOS Transistor (BSIM4 Model)
M2 out in vdd vdd PMOS L='tplv' W='tpwv'
.model PMOS pmos level=54
+ toxe=tpotv                * PMOS transistor oxide thickness variation
+ ...                       * Additional PMOS BSIM4 parameters as needed

* Load Capacitance
Cload out 0 1p

* Simulation Control
.tran 1n 100n
.end
